*This is a sample input deck for SCAPP
v1 1 0 DC 0 AC 1

r1 1 2 1
c1 2 0 1
r4 2 3 1
c2 3 0 1
l5 3 4 1
c3 4 0 1
r6 4 5 1
c6 5 0 1
.AC DEC 1 1 10
.PRINT ac vdb(5)
.end
