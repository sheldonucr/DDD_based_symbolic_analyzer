CMOS OPAMP
*
VDD 1 0 DC 5 
*VAP 34 99 PULSE( 0.0 0.5 0 1e-9 1e-9 50e-9 100e-9)
*VAP 34 99 AC 1
*Vin 99 0 dc 2.5
VIN 34 0 DC 2.5 AC 1
*
*
* ANALOG INOUT
*
*BASIC CIRCUIT

M65	0 0 7 1 PCH W=4.5u L=40u
M64	7 7 1 1 PCH W=71u L=10u
M63	5 7 1 1 PCH W=69u L=10u
M62	5 5 9 0 NCH W=35u L=10u
M61	9 9 0 0 NCH W=12u L=10u
*
* Differentail amplifier stage
*
M10 36 33 32 1 PCH W=11u L=2u AD=24p AS=24p
M20 3 34 32 1 PCH W=11u L=2u AD=24p AS=24p
M30 36 36 0 0 NCH w=6u l=3u AD=136p as=136p
M40 3 36 0 0 NCH W=6u L=3u AD=136p AS=136p
M50 32 7 1 1 PCH W=14u L=2u AD=24p AS=24p

*
* Folded cascode stage with compensation
*
M2 6 7 1 1 PCH W=80u L=2u AD=24p AS =24p
M3 6 5 4 0 NCH w=24u L=2u AD=136p AS=136p
M4 4 3 0 0 NCH w=46u L=2u AD=136p AS=136p
M80 11 5 3 0 NCH w=4u L=3u 
CC 6 11 .22pf

* Common drain output stage
M7 1 6 12 12 NCH W=100u L=2u AD=136p AS=136p
M8 12 9 0 0 NCH W=63u L=2u AD=136p AS=136p

* load
CL 12 0 10pf

* feedback
RF 12 33 100
*
* MOSFET PROCESS MODEL
*
.MODEL NCH NMOS LEVEL=2  VTO=0.9 KP=50E-6 GAMMA=0.30 PHI=0.70
+ CGSO=1.76E-10 CGDO=1.76E-10 CJ=0.7E-4 MJ=0.5 CJSW=3.9E-10 MJSW=0.33 JS=1E-3
+ TOX=42.5N NFS=1E11 LD=0 UCRIT=1E4
+ LAMBDA=0.019

.MODEL N NMOS LEVEL=2 CGSO=2.89E-10 VTO=0.71 GAMMA=0.29
+ CGDO=2.89E-10 CJ=3.74E-4 TOX=225E-10 NSUB=3.5E16
+ UO=411 LAMBDA=0.02

.MODEL PCH PMOS LEVEL=2 VTO=-0.9 KP=17E-6 GAMMA=0.50 PHI=0.69
+ CGSO=2.8E-10 CGDO=2.8E-10 CJ=3.3E-4 MJ=0.5 CJSW=4.4E-10 MJSW=0.33 JS=1E-3
+ TOX=42.5N LD=0 UCRIT=1E4 NFS=1E11
+ LAMBDA=0.005

.MODEL P PMOS LEVEL=2 VTO=-0.76 GAMMA=0.6 CGSO=3.35E-10
+CGDO=3.35E-10 CJ=4.75E-4 MJ=0.4 TOX=225E-10 NSUB=1.6E16 
+ XJ=0.2E-6 UO=139 LAMBDA=0.02

*
*
*
*.OP
*.OPTIONS ACCT ITL1=300
.AC DEC 10 1 100M 
.PRINT VDB(12)
.END
