*
r1 1 2 10k
r2 2 0 5k
r3 2 3 5k
r4 3 0 10k
r5 3 4 5k
r6 4 0 5k
In 1 0 DC 0 AC 1
.AC DEC 100 100 1000
.print ac vdb(4)
.end

