*This is a RC ladder tree 
*#(top level)total nodes (DDD): 301
*#nodes (DDD): 98
*#paths (DDD): 142400
*#nodes (DDD): 225
*#paths (DDD): 3.02514e+10


R1 1 0 1k
c2 1 2 1k
R3 2 0 1k
r4 2 3 1k
c5 3 0 1k
c6 3 4 1k
R7 4 0 1k
R8 4 5 1k
c9 5 0 1k
R10 5 6 1k
c11 6 0 1k
R12 6 7 1k
c13 7 0 1k
c14 7 8 1k
c15 8 0 1k
R16 8 9 1k
c17 9 0 1k
R18 9 10 1k
c19 10 0 1k
R20 10 11 1k

R21 11 0 1k
c22 11 12 1k
R23 12 0 1k
R24 12 13 1k
c25 13 0 1k
R26 13 14 1k
c27 14 0 1k
R28 14 15 1k
c29 15 0 1k

R30 11 16 1k
c31 16 0 1k
R32 16 17 1k
c33 17 0 1k
r34 17 18 1k
c35 18 0 1k
r36 18 19 1k
R37 19 0 1k
r38 19 20 1k
c39 20 0 1k

c40 11 21 1k
R41 21 0 1k
r42 21 22 1k
r43 22 0 1k
c44 22 23 1k
R45 23 0 1k
c46 23 24 1k
R47 24 0 1k
c48 24 25 1k
R49 25 0 1k
c50 25 26 1k
R51 26 0 1k
c52 26 27 1k
R53 27 0 1k
c54 27 28 1k
R55 28 0 1k
c56 28 29 1k
R57 29 0 1k
c58 29 30 1k
R59 30 0 1k

c60 11 31 1k
R61 31 0 1k
c62 31 32 1k
R63 32 0 1k
r64 32 33 1k
c65 33 0 1k
R66 33 34 1k
c67 34 0 1k
c68 34 35 1k
R69 35 0 1k
c70 35 36 1k
R71 36 0 1k
c72 36 37 1k
R73 37 0 1k
c74 37 38 1k
R75 38 0 1k
c76 38 39 1k
R77 39 0 1k
c78 39 40 1k
R79 40 0 1k


R80 40 41 1k
c81 41 0 1k
R82 41 42 1k
c83 42 0 1k
r84 42 43 1k
r85 43 0 1k
c86 43 44 1k
R87 44 0 1k

R100 40 51 1k
c101 51 0 1k
R102 51 52 1k
c103 52 0 1k
c104 52 53 1k
R105 53 0 1k
c106 53 54 1k
R107 54 0 1k

R120 40 61 1k
c121 61 0 1k
R122 61 62 1k
c123 62 0 1k
c124 62 63 1k
R125 63 0 1k
c126 63 64 1k
R127 64 0 1k
c128 64 65 1k
R129 65 0 1k

g1 1 0 44 0 0
vin 1 0 dc 0 ac 1
.ac dec 1000 1 10
.plot vdb(44)
.end
