*This is a sample input deck for SCAPP
v1 10 0 DC 0 AC 1
r1 10 1 0.5k
c1 1 0 2u
r2 1 2 1k
c2 2 0 1u
r3 2 3 1k
c3 3 0 1u
.AC DEC 100 100 1000 
.print ac v(3)
.end
