* This file coming from the Starzyk's bandpass example
* modified in May 26, 1998
r1 1 2 1 
r2 12 8 1 
r3 2 0 1
rr 2 3 1
r4 8 3 1
r5 3 4 1
r6 4 5 1
c6 4 5 1
r7 5 6 1
c8 6 7 1
r9 7 8 1
r10 5 9 1 
r11 19 15 1 
r12 9 0 1
rr1 9 10 1
r13 10 15 1
r14 10 11 1
r15 11 12 1
c15 11 12 1
r16 12 13 1
c17 13 14 1
r18 14 15 1
r19 12 16 1
rr2 16 17 1
r20 22 26 1
r21 16 0 1
r22 22 17 1
r23 17 18 1
r24 18 19 1
c24 18 19 1
r25 19 20 1
c26 20 21 1
r27 21 22 1
r28 19 23 1
r29 29 30 1
r30 23 0 1
r31 24 29 1
r32 24 25 1
r33 25 26 1
c33 25 26 1
r34 26 27 1
c35 27 28 1
r36 28 29 1
r37 26 31 1
r38 32 0 1
r39 31 0 1
r40 32 30 1

r41 23 22 1
c42 23 32 1
rr3 15 16 1
l43 11 12 1
*l44 22 26 1
r49 17 28 1
c46 16 21 1

*r45 24 2 1
*c43 21 26 1
*l47 10 9 1
*l42 20 21 1
g11 1 0 32 0 0.0

v1 1 0 DC 0 AC 1 
.AC DEC 2  1 100meg 
.PRINT ac vdb(32) vdb(33) vdb(23)
.end
