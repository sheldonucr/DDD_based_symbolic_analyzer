*************************************
* DETAILED CIRCUIT FROM BOYLE PAPER *
*************************************
.SUBCKT UA741  1 2 24 27 26
* NODES: IN+ IN- OUT VCC VEE
R1 10 26 1K
R2 9 26 50K
R3 11 26 1K
R4 12 26 3K
R5 15 17 39K
R6 23 24 50
R7 24 25 25
R8 18 26 100
R9 14 26 50K
R10 21 20 40K
R11 13 26 50K
COMP 22 8 30PF
Q1 3 1 4 BNP1
Q2 3 2 5 BNP1
Q3 7 6 4 BPN1
Q4 8 6 5 BPN1
Q5 7 9 10 BNP1
Q6 8 9 11 BNP1
Q7 27 7 9 BNP1
Q8 3 3 27 BPN1
Q9 6 3 27 BPN1
Q10 6 15 12 BNP1
Q11 15 15 26 BNP1
Q12 17 17 27 BPN1
Q13A 28 17 27 BPN3
Q13B 22 17 27 BPN4
Q14 27 28 23 BNP2
Q15 28 23 24 BNP1
Q16 27 8 14 BNP1
Q17 22 14 18 BNP1
Q18 28 21 20 BNP1
Q19 28 28 21 BNP1
Q20 26 20 25 BPN2
Q21 13 25 24 BPN1
Q22 8 13 26 BNP1
Q23A 26 22 20 BPN5
Q23B 26 22 8 BPN6
Q24 13 13 26 BNP1
*
.MODEL BNP1 NPN BF=209 BR=2.5 RB=670 RC=300 CCS=1.417P TF=1.15N TR=405N
+ CJE=0.65P CJC=0.36P IS=1.26E-15 VA=178.6 IK=1.611M NE=2 PE=0.6
+ ME=0.33 PC=0.45 MC=0.33
.MODEL BNP2 NPN BF=400 BR=6.1 RB=185 RC=15 CCS=3.455P TF=0.76N TR=243N
+ CJE=2.80P CJC=1.55P IS=0.395E-15 VA=267 IK=10M NE=2 PE=0.6
+ ME=0.33 PC=0.45 MC=0.33
.MODEL BPN1 PNP BF=75 BR=3.8 RB=500 RC=150 CCS=2.259P TF=27.4N TR=2540N
+ CJE=0.10P CJC=1.05P IS=3.15E-15 VA=55.11 IK=270U NE=2 PE=0.45
+ ME=0.33 PC=0.45 MC=0.33
.MODEL BPN2 PNP BF=117 BR=4.8 RB=80 RC=156 TF=27.4N TR=2540N
+ CJE=4.05P CJC=2.80P IS=17.6E-15 VA=57.94 IK=590.7U NE=2 PE=0.6
+ ME=0.25 PC=0.6 MC=0.25
.MODEL BPN3 PNP BF=13.8 BR=1.4 RB=100 RC=80 CCS=2.126P TF=27.4N TR=55N
+ CJE=0.10P CJC=0.3P IS=2.25E-15 VA=83.55 IK=5M NE=2 PE=0.45
+ ME=0.33 PC=0.45 MC=0.33
.MODEL BPN4 PNP BF=14.8 BR=1.5 RB=160 RC=120 CCS=2.126P TF=27.4N TR=220N
+ CJE=0.10P CJC=0.90P IS=2.25E-15 VA=83.55 IK=171.8U NE=2 PE=0.45
+ ME=0.33 PC=0.45 MC=0.33
.MODEL BPN5 PNP BF=80 BR=1.5 RB=1100 RC=170 TF=26.5N TR=9550N
+ CJE=0.10P CJC=2.40P IS=0.79E-15 VA=79.45 IK=80.55U NE=2 PE=0.6
+ ME=0.25 PC=0.6 MC=0.25
.MODEL BPN6 PNP BF=19 BR=1.0 RB=650 RC=100 TF=26.5N TR=2120N
+ CJE=1.90P CJC=2.40P IS=0.63E-17 VA=167.1 IK=80.55U NE=2 PE=0.6
+ ME=0.25 PC=0.6 MC=0.25
*
.ENDS UA741
*********************
* UA741 MACRO-MODEL *
*********************
.SUBCKT UA741MAC 3 2 6 7 4
* NODES: IN+ IN- OUT VCC VEE
Q1 8 2 10 QMOD1
Q2 9 3 11 QMOD2
RC1 7 8 4352
RC2 7 9  4352
RE1 1 10 2391.9
RE2 1 11 2391.9
RE 1 0 7.27MEG
CE 1 0 7.5P
IEE 1 4 27.512U
C1 8 9 4.5288P
RP 7 4 15.363K
GCM 0 12 1 0 1.1516N
GA 12 0 8 9 229.774U
R2 12 0 100K
C2 12 13 30P
GB 13 0 12 0 37.0978
R02 13 0 489.2
R01 13 6 76.8
D1 13 14 DMOD1
D2 14 13 DMOD1
EC 0 14 6 0 1
*GC 0 14 6 0 5034.3
RC 14 0 0.1986M
D3 6 15 DMOD3
D4 16 6 DMOD3
VC 7 15 1.6042
VE 16 4 3.1042
*
.MODEL QMOD1 NPN IS=8E-16 BF=52.6726
.MODEL QMOD2 NPN IS=8.0925E-16 BF=52.7926
.MODEL DMOD1 D IS=3.8218E-32
.MODEL DMOD3 D IS=8E-16
.ENDS
*UA741 FREQUENCY RESPONSE
*
* MACRO MODEL
X1 1 0 3 4 5 UA741MAC
* FULL MODEL
X2 2 0 6 4 5 UA741
*
VIN1 1 0 DC -.2765M AC 1
VIN2 2 0 DC -.2834M AC 1
VCC 4 0 15
VEE 5 0 -15
*
*
.TF V(3) VIN1
.TF V(6) VIN2
.AC DEC 10 .1 1G
.END

