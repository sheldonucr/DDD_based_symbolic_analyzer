*This is the example used in our paper. 5/24/02
r1 1 0 5k
c1 1 0 2u
r2 1 2 2k
c2 2 0 4u
r3 2 3 3k
c3 3 0 8u
I1 1 0 DC 10mA 
.AC DEC 5 100 1000 
.print ac v(3)
.end
