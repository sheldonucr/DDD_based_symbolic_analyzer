*
r1 1 2 10k
c1 1 0 10u
c2 2 0 20u
in 1 0 DC 0 AC 1
.AC DEC 100 100 1e6
.print ac vdb(2)
.end

