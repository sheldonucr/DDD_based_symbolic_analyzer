*single stage amplifer
*mxxx d g s b
M2A   3 2 0 0 N W=100U L=20.3U AD=99P   AS=99P   PD=40U   PS=40U
RL 3 0 5k
RS 1 2 100k
CL 1 2 10p

VIN 1 0 DC 3 AC 1 
VDD 4 0 DC 5
I1 4 3 DC 10m

.MODEL N NMOS LEVEL=2  VTO=0.9 KP=50E-6 GAMMA=0.30 PHI=0.70
+ CGSO=1.76E-10 CGDO=1.76E-10 CJ=0.7E-4 MJ=0.5 CJSW=3.9E-10 MJSW=0.33 JS=1E-3
+ TOX=42.5N NFS=1E11 LD=0 UCRIT=1E4
+ LAMBDA=0.019

*.OP
.AC DEC 10 1 100MEG
.END
