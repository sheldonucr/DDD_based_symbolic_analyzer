*This is a sample input deck for SCAPP
v1 1 0 DC 0 AC 1
r1 1 2 5meg
l1 2 0 20m
.AC DEC 100 100 1000 
.print ac vdb(2)
.end
