*This is a sample input deck for SCAPP
v1 1 0 DC 0 AC 1
r1 1 2 5k
c1 2 0 2u
r2 2 3 2k
c2 3 0 4u
r3 3 4 3k
c3 4 0 8u
.AC DEC 5 100 1000 
.print ac v(4)
.end
