*This is is an exmaple
R1 1 3 1k
c2 3 0 1pf
cc3 1 2 1pf
R4 2 4 1k
c5 4 0 1pf
R6 3 5 1k
c7 5 0 1pf
cc8 3 4 1pf
R9 4 6 1k
c10 6 0 1pf
R11 5 7 1k
c12 7 0 1pf
cc13 5 6 1pf
R14 6 8 1k
c15 8 0 1pf
R16 7 9 1k
c17 9 0 1pf
cc18 7 8 1pf
R19 8 10 1k
c20 10 0 1pf
R21 9 11 1k
c22 11 0 1pf
cc23 9 10 1pf
R24 10 12 1k
c25 12 0 1pf
R26 11 13 1k
c27 13 0 1pf
cc28 11 12 1pf
R29 12 14 1k
c30 14 0 1pf
R31 13 15 1k
c32 15 0 1pf
cc33 13 14 1pf
R34 14 16 1k
c35 16 0 1pf
R36 15 17 1k
c37 17 0 1pf
cc38 15 16 1pf
vin 2 0 dc 0 ac 1
.ac dec 10 10  10000
.plot vdb(16)
.end
